// tb_uart_top.sv

`default_nettype none

module tb_uart_top;

initial begin
  run_test();
end

endmodule
